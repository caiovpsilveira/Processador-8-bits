library verilog;
use verilog.vl_types.all;
entity simulacao_processador is
end simulacao_processador;
